-- font_ufm.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity font_ufm is
	port (
		addr       : in  std_logic_vector(8 downto 0)  := (others => '0'); --       addr.addr
		data_valid : out std_logic;                                        -- data_valid.data_valid
		dataout    : out std_logic_vector(15 downto 0);                    --    dataout.dataout
		nbusy      : out std_logic;                                        --      nbusy.nbusy
		nread      : in  std_logic                     := '0'              --      nread.nread
	);
end entity font_ufm;

architecture rtl of font_ufm is
	component font_ufm_ufm_parallel_0 is
		port (
			addr       : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- addr
			nread      : in  std_logic                     := 'X';             -- nread
			dataout    : out std_logic_vector(15 downto 0);                    -- dataout
			nbusy      : out std_logic;                                        -- nbusy
			data_valid : out std_logic                                         -- data_valid
		);
	end component font_ufm_ufm_parallel_0;

begin

	ufm_parallel_0 : component font_ufm_ufm_parallel_0
		port map (
			addr       => addr,       --       addr.addr
			nread      => nread,      --      nread.nread
			dataout    => dataout,    --    dataout.dataout
			nbusy      => nbusy,      --      nbusy.nbusy
			data_valid => data_valid  -- data_valid.data_valid
		);

end architecture rtl; -- of font_ufm
